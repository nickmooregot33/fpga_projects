module counter();


endmodule
