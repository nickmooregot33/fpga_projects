module test_tb;

test_top dut();


endmodule
